module clk_div (
	input wire i_ref_clk, i_rst_n, i_clk_en,
	input wire [3:0] i_div_ratio,
	output reg o_div_clk
	);

reg [2:0] counter;
reg count_up_done, count_dn_done;

wire [2:0] up_counts;
wire [3:0] dn_counts;

assign up_counts = i_div_ratio[3:1];
assign dn_counts = (i_div_ratio[0] == 1'b0 )? up_counts : up_counts+1;

always @(posedge i_ref_clk or negedge i_rst_n) begin
	
	if (! i_rst_n) begin
		counter<='b0;
        count_up_done<=1'b0;
        count_dn_done<=1'b0;
        o_div_clk<=1'b0;
	end
	else if (i_clk_en & (i_div_ratio != 'b0 & i_div_ratio != 'b1) & !count_up_done) begin
		o_div_clk<=1'b1;
		counter<=counter+1;
		if(counter== up_counts-1) begin
			counter<='b0;
			count_up_done<=1'b1;
			count_dn_done<=1'b0;
		end
	end
	else if (i_clk_en & (i_div_ratio != 'b0 & i_div_ratio != 'b1) & !count_dn_done) begin
        o_div_clk<=1'b0;
        counter<=counter+1;
		if(counter== dn_counts-1) begin
			counter<='b0;
			count_up_done<=1'b0;
			count_dn_done<=1'b1;
		end
	end
	else begin
	    o_div_clk<=1'b0;
		counter<='b0;
        count_up_done<=1'b0;
        count_dn_done<=1'b0;
	end
end


endmodule